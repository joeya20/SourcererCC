begin
        reg_rdata_next[31:0] = reg2hw.key_share0[0].q;
      end