assign wipe_secret_we = addr_hit[8] & reg_we & reg_error;
