begin
  if (counter_done) state_d = Done;
end
